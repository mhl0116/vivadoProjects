
// file: ibert_ultrascale_gth_0.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_ultrascale_gth_0
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_ultrascale_gth_0
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 1
`define C_GTH_REFCLKS_USED 1
module example_ibert_ultrascale_gth_0
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txn_o,
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txp_o,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]    	gth_rxn_i,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]   	gth_rxp_i,
  input                           	gth_sysclkp_i,
  input                           	gth_sysclkn_i,
  output                            sel_si750_clk_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0n_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1n_i,
  output reg [1:0]                          gpio_led
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;        	
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i; 
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                        gth_sysclk_i;


  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE3 u_buf_gth_q3_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[0]),
        .IB           (gth_refclk0n_i[0])
      );
    IBUFDS_GTE3 u_buf_gth_q3_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[0]),
        .IB           (gth_refclk1n_i[0])
      );

  //
  wire clk_out40;
    
  clockManager clockManager_i
   (
    // Clock out ports
    .clk_out1(clk_out40),     // output clk_out1
    // Clock in ports
    .clk_in1(gth_sysclk_i)
    );      // input clk_in300
    
  reg div_temp;
  wire reset;
  reg[15:0] cnt;
  
  always @ (posedge clk_out40) begin
    
    if (reset) begin
        cnt <= 16'b0;
    end else if (cnt == 16'hFFFF) begin
        div_temp <= !div_temp;
        cnt <= cnt + 1'b1; 
    end else begin
    cnt <= cnt + 1'b1;
    end
    
    gpio_led[0] <= div_temp;
    
  end
    
  wire [31:0] ila_data; 
  wire [7:0] ila_trigger; 
  
  assign ila_data[0] = reset;
  assign ila_data[1] = div_temp;
  assign ila_data[17:2] = cnt;
  
  assign ila_trigger[1] = div_temp;
  assign ila_trigger[0] = reset;
  
  ila_0 ila_i (
	.clk(clk_out40), // input wire clk

	.probe1(ila_trigger), // input wire [7:0]  probe0  
	.probe0(ila_data) // input wire [31:0]  probe1
  );
  
  
  vio_0 vio_i (
    .clk (clk_out40)
    ,.probe_out0 (reset)
  );
    
  assign sel_si750_clk_i = 1'b0;
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = 1'b0;
  assign gth_qrefclk1_i[0] = 1'b0;
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = 1'b0;
  assign gth_qrefclk10_i[0] = 1'b0;
  assign gth_qrefclk01_i[0] = 1'b0;
  assign gth_qrefclk11_i[0] = 1'b0;
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;
  assign gth_qsouthrefclk00_i[0] = gth_refclk0_i[0];
  assign gth_qsouthrefclk10_i[0] = 1'b0;
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0;
 
  //
  // Sysclock IBUFDS instantiation
  //
  IBUFGDS 
   #(.DIFF_TERM("FALSE"))
   u_ibufgds
    (
      .I(gth_sysclkp_i),
      .IB(gth_sysclkn_i),
      .O(gth_sysclk_i)
    );


  //
  // IBERT core instantiation
  //
  ibert_ultrascale_gth_0 u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(gth_sysclk_i),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

endmodule
